package alu_type is
	type TYPE_OP is (ADD, SUB, BITAND, BITOR);
	--type TYPE_OP is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, FUNCRL, FUNCRR);
end alu_type;
