package CONSTANTS is
   constant IVDELAY : time := 0.1 ns;
   constant NDDELAY : time := 0.2 ns;
   constant NDDELAYRISE : time := 0.6 ns;
   constant NDDELAYFALL : time := 0.4 ns;
   constant NRDELAY : time := 0.2 ns;
   constant DRCAS : time := 0 ns;
   constant DRCAC : time := 0 ns;
   constant numBit : integer := 32;	
   constant tp_mux : time := 0.5 ns; 
   constant NBIT_PER_BLOCK : integer := 4;
   --constant NBLOCKS	: integer := 8;
   constant NBIT: integer := 32;
end CONSTANTS;
