111101100000101--ADD
101000100000101--ADDI
111101100000101--AND
101000100000101--ANDI
101000101100100--BEQZ
101000101100100--BNEZ
101000110000001--J
101010110000001--JAL
001000100000101--LW
001000100000100--NOP
111101100000101--OR
101000100000101--ORI
000000000000000--SGE
000000000000000--SGEI
000000000000000--SLE
000000000000000--SLEI
000000000000000--SLL
000000000000000--SLLI
000000000000000--SNE
000000000000000--SNEI
000000000000000--SRL
000000000000000--SRLI
111101100000101--SUB
101000100000101--SUBI
000000000000000--SW
111101100000101--XOR
101000100000101--XORI





--RF1,	RF2,	EN1,	I0_R1_SEL,	JAL_SEL,	I0_R1_S2,		EN2,	ISJUMP,	ISBRANCH,	BEQZ,	RM,	WM,	EN3,	S3_1M_0ALU,	WF1
--0,	1,  	2,		3,			4,			5,				6,		7,		8,			9,		10,	11,	12,		13, 		14
